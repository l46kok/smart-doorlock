CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
680 0 30 200 10
176 80 1678 989
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
31
5 SIP4~
219 927 20 0 4 9
0 5 4 3 2
0
0 0 608 90
4 CONN
9 2 37 10
2 J9
-10 -19 4 -11
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 J
7849 0 0
2
42690.7 0
0
9 Schottky~
219 462 44 0 2 5
0 8 16
0
0 0 832 0
8 SCHOTTKY
-27 -18 29 -10
2 D2
-6 -28 8 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6343 0 0
2
5.89777e-315 0
0
9 Schottky~
219 378 177 0 2 5
0 11 9
0
0 0 832 90
8 SCHOTTKY
12 -1 68 7
2 D1
33 -11 47 -3
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7376 0 0
2
5.89777e-315 0
0
9 Schottky~
219 252 138 0 2 5
0 10 9
0
0 0 832 0
8 SCHOTTKY
-27 -18 29 -10
2 D4
-6 -28 8 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9156 0 0
2
5.89777e-315 0
0
10 N-EMOS 3T~
219 427 65 0 3 7
0 8 7 6
0
0 0 832 0
11 IRLB8721PbF
8 0 85 8
2 Q1
28 -10 42 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
4 SIP3
7

0 2 1 3 2 1 3 0
77 0 0 0 1 1 0 0
1 Q
5776 0 0
2
5.89777e-315 0
0
5 SIP2~
219 396 125 0 2 5
0 9 16
0
0 0 1632 90
4 CONN
9 2 37 10
2 J1
-15 -19 -1 -11
12 Power Switch
-71 -28 13 -20
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
7207 0 0
2
42690.7 0
0
5 SIP3~
219 206 149 0 3 7
0 18 6 10
0
0 0 1632 180
4 CONN
-13 -25 15 -17
2 J3
-10 -26 4 -18
9 9V (Wall)
-31 -35 32 -27
0
0
0
0
8 PCBPower
7

0 3 1 2 3 1 2 0
0 0 0 512 1 1 0 0
1 J
4459 0 0
2
42690.7 1
0
5 SIP3~
219 331 257 0 3 7
0 19 6 11
0
0 0 1632 180
4 CONN
-13 -25 15 -17
2 J8
-12 -25 2 -17
11 7.2V (Batt)
-43 -34 34 -26
0
0
0
0
8 PCBPower
7

0 3 1 2 3 1 2 0
0 0 0 512 1 1 0 0
1 J
3760 0 0
2
42690.7 2
0
5 SIP6~
219 968 45 0 6 13
0 12 5 4 3 2 6
0
0 0 1632 0
4 CONN
9 2 37 10
2 J7
-7 -38 7 -30
20 Keypad / Buzzer GPIO
-17 33 123 41
0
0
0
0
4 SIP6
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
0 0 0 0 1 0 0 0
1 J
754 0 0
2
5.89777e-315 0
0
5 SIP2~
219 707 56 0 2 5
0 14 13
0
0 0 1632 0
4 CONN
9 2 37 10
2 J6
-7 -20 7 -12
11 Buzzer (5V)
-31 -30 46 -22
0
0
0
0
6 RAD0.3
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 J
9767 0 0
2
5.89777e-315 5.26354e-315
0
10 N-EMOS 3T~
219 680 93 0 3 7
0 14 12 6
0
0 0 832 0
6 VN2106
18 0 60 8
2 Q2
32 -10 46 -2
0
0
17 %D %1 %2 %3 %3 %M
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
77 0 0 256 1 0 0 0
1 Q
7978 0 0
2
5.89777e-315 5.30499e-315
0
5 SIP3~
219 212 67 0 3 7
0 17 8 16
0
0 0 1632 180
4 CONN
-13 -25 15 -17
2 J4
-10 -26 4 -18
19 Solenoid Power/GPIO
-28 16 105 24
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
3142 0 0
2
5.89777e-315 5.32571e-315
0
10 Polar Cap~
219 858 192 0 2 5
0 15 6
0
0 0 832 270
5 100uF
2 6 37 14
2 C6
14 -6 28 2
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3284 0 0
2
5.89777e-315 5.34643e-315
0
10 Polar Cap~
219 284 189 0 2 5
0 9 6
0
0 0 832 270
5 470uF
5 8 40 16
2 C1
10 -4 24 4
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
659 0 0
2
5.89777e-315 5.3568e-315
0
5 SIP4~
219 924 206 0 4 9
0 15 15 6 6
0
0 0 1632 0
4 CONN
9 2 37 10
2 J2
-7 -29 7 -21
20 MCU/NFC Power (3.3V)
-25 -38 115 -30
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 J
3800 0 0
2
5.89777e-315 5.38788e-315
0
5 SIP4~
219 676 204 0 4 9
0 13 13 6 6
0
0 0 1632 0
4 CONN
9 2 37 10
2 J5
-7 -29 7 -21
21 LCD/Keypad Power (5V)
-59 28 88 36
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
1 J
6792 0 0
2
5.89777e-315 5.40342e-315
0
10 Polar Cap~
219 820 160 0 2 5
0 15 6
0
0 0 832 270
4 22uF
9 8 37 16
2 C5
10 -4 24 4
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3701 0 0
2
5.89777e-315 5.4086e-315
0
10 Polar Cap~
219 714 169 0 2 5
0 13 6
0
0 0 832 270
4 10uF
9 8 37 16
2 C4
10 -4 24 4
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6316 0 0
2
5.89777e-315 5.41378e-315
0
11 Regulator3~
219 759 148 0 3 7
0 13 6 15
0
0 0 4928 0
13 LT1805 CT-3.3
-46 -28 45 -20
2 U3
-7 -38 7 -30
0
0
14 %D %1 %2 %3 %S
0
0
4 SIP3
7

0 3 1 2 3 1 2 0
88 0 0 0 1 1 0 0
1 U
8734 0 0
2
5.89777e-315 5.41896e-315
0
10 Polar Cap~
219 614 166 0 2 5
0 13 6
0
0 0 832 270
5 0.1uF
4 9 39 17
2 C3
10 -4 24 4
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7988 0 0
2
42690.7 3
0
10 Polar Cap~
219 501 164 0 2 5
0 16 6
0
0 0 832 270
6 0.33uF
2 8 44 16
2 C2
10 -4 24 4
0
0
11 %D %1 %2 %V
0
0
4 SIP2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3217 0 0
2
42690.7 4
0
11 Regulator3~
219 561 147 0 3 7
0 16 6 13
0
0 0 4928 0
8 OKI-78SR
-28 -28 28 -20
2 U2
-7 -38 7 -30
0
0
14 %D %1 %2 %3 %S
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
88 0 0 0 1 0 0 0
1 U
3965 0 0
2
42690.7 5
0
7 Ground~
168 451 298 0 1 3
0 20
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
8239 0 0
2
42690.7 6
0
9 Resistor~
219 411 103 0 2 5
0 6 7
0
0 0 864 90
4 100k
2 0 30 8
2 R8
6 -10 20 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
828 0 0
2
5.89777e-315 0
0
9 Resistor~
219 610 99 0 2 5
0 6 12
0
0 0 864 90
4 100k
4 0 32 8
2 R7
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6187 0 0
2
5.89777e-315 5.42414e-315
0
9 Resistor~
219 829 32 0 2 5
0 15 5
0
0 0 864 0
3 10k
-10 -14 11 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7107 0 0
2
5.89777e-315 5.42933e-315
0
9 Resistor~
219 829 113 0 2 5
0 15 2
0
0 0 864 0
3 10k
-11 -12 10 -4
2 R5
-7 -21 7 -13
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6433 0 0
2
5.89777e-315 5.43192e-315
0
9 Resistor~
219 828 87 0 2 5
0 15 3
0
0 0 864 0
3 10k
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8559 0 0
2
5.89777e-315 5.43451e-315
0
9 Resistor~
219 829 57 0 2 5
0 15 4
0
0 0 864 0
3 10k
-11 -11 10 -3
2 R3
-8 -20 6 -12
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3674 0 0
2
5.89777e-315 5.4371e-315
0
9 Resistor~
219 366 74 0 2 5
0 17 7
0
0 0 864 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5697 0 0
2
5.89777e-315 5.43969e-315
0
9 Resistor~
219 333 179 0 2 5
0 11 9
0
0 0 864 90
2 1k
6 -5 20 3
2 R1
5 -14 19 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3805 0 0
2
42690.7 7
0
61
4 0 2 0 0 4096 0 1 0 0 32 2
938 29
938 59
3 0 3 0 0 4096 0 1 0 0 33 2
929 29
929 50
2 0 4 0 0 4096 0 1 0 0 34 2
920 29
920 41
1 0 5 0 0 12288 0 1 0 0 35 4
911 29
911 28
911 28
911 32
1 0 6 0 0 8192 0 24 0 0 21 3
411 121
411 125
433 125
0 2 7 0 0 4096 0 0 24 51 0 3
403 74
403 85
411 85
1 0 8 0 0 4096 0 2 0 0 30 2
451 44
433 44
2 0 9 0 0 4096 0 3 0 0 48 2
379 164
379 138
1 3 10 0 0 4224 0 4 7 0 0 2
241 138
213 138
0 2 9 0 0 0 0 0 4 53 0 2
271 138
264 138
4 0 6 0 0 4096 0 15 0 0 59 2
912 220
857 220
2 0 6 0 0 8192 0 17 0 0 14 3
819 167
819 193
759 193
2 0 6 0 0 0 0 18 0 0 14 2
713 176
759 176
2 0 6 0 0 4096 0 19 0 0 59 2
759 172
759 283
0 0 6 0 0 4096 0 0 0 25 59 2
686 123
686 283
4 0 6 0 0 0 0 16 0 0 20 2
664 218
561 218
3 0 6 0 0 0 0 16 0 0 20 2
664 209
561 209
2 0 6 0 0 0 0 20 0 0 20 3
613 173
613 184
561 184
2 0 6 0 0 0 0 21 0 0 20 3
500 171
500 194
561 194
2 0 6 0 0 0 0 22 0 0 59 2
561 171
561 283
3 0 6 0 0 4096 0 5 0 0 59 2
433 83
433 283
2 0 6 0 0 0 0 14 0 0 59 2
283 196
283 283
0 2 6 0 0 0 0 0 8 59 0 3
356 283
356 255
338 255
0 3 11 0 0 4096 0 0 8 60 0 3
356 214
356 246
338 246
1 3 6 0 0 0 0 25 11 0 0 4
610 117
610 123
686 123
686 111
0 2 12 0 0 4096 0 0 25 29 0 3
654 75
610 75
610 81
2 0 13 0 0 4096 0 10 0 0 57 2
695 61
695 139
1 1 14 0 0 8320 0 10 11 0 0 3
695 52
686 52
686 75
1 2 12 0 0 8320 0 9 11 0 0 5
956 23
956 5
654 5
654 102
662 102
1 2 8 0 0 8320 0 5 12 0 0 5
433 47
433 34
227 34
227 65
219 65
0 1 13 0 0 0 0 0 19 57 0 2
713 139
731 139
5 2 2 0 0 4224 0 9 27 0 0 4
956 59
875 59
875 113
847 113
4 2 3 0 0 4224 0 9 28 0 0 4
956 50
859 50
859 87
846 87
3 2 4 0 0 4224 0 9 29 0 0 4
956 41
855 41
855 57
847 57
2 2 5 0 0 4224 0 9 26 0 0 2
956 32
847 32
6 0 6 0 0 0 0 9 0 0 59 6
956 68
914 68
914 118
1037 118
1037 283
857 283
1 0 15 0 0 4096 0 28 0 0 41 2
810 87
805 87
1 0 15 0 0 4096 0 27 0 0 41 2
811 113
805 113
1 0 15 0 0 0 0 29 0 0 41 2
811 57
805 57
1 0 15 0 0 0 0 26 0 0 41 3
811 32
805 32
805 31
0 0 15 0 0 4224 0 0 0 56 40 2
805 139
805 31
1 0 13 0 0 0 0 16 0 0 52 2
664 191
654 191
1 3 13 0 0 0 0 20 22 0 0 3
613 156
613 138
589 138
3 0 6 0 0 0 0 15 0 0 59 2
912 211
857 211
1 0 15 0 0 0 0 13 0 0 56 3
857 182
857 178
893 178
2 0 15 0 0 0 0 15 0 0 56 3
912 202
893 202
893 193
0 1 16 0 0 4096 0 0 22 58 0 2
500 138
533 138
0 1 9 0 0 4224 0 0 6 61 0 3
333 138
389 138
389 134
1 0 15 0 0 0 0 17 0 0 56 2
819 150
819 139
1 1 17 0 0 4224 0 30 12 0 0 2
348 74
219 74
2 2 7 0 0 4224 0 5 30 0 0 2
409 74
384 74
2 0 13 0 0 0 0 16 0 0 57 3
664 200
654 200
654 139
0 1 9 0 0 0 0 0 14 0 0 3
268 138
283 138
283 179
0 2 16 0 0 8192 0 0 6 55 0 4
488 56
488 138
398 138
398 134
3 2 16 0 0 12416 0 12 2 0 0 8
219 56
224 56
224 25
503 25
503 56
481 56
481 44
474 44
3 1 15 0 0 0 0 19 15 0 0 4
787 139
893 139
893 193
912 193
1 0 13 0 0 8320 0 18 0 0 43 3
713 159
713 139
613 139
1 0 16 0 0 0 0 21 0 0 54 3
500 154
500 138
488 138
2 2 6 0 0 12416 0 7 13 0 0 5
213 147
225 147
225 283
857 283
857 199
1 1 11 0 0 8320 0 3 31 0 0 4
379 187
379 214
333 214
333 197
2 0 9 0 0 0 0 31 0 0 53 3
333 161
333 138
283 138
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
429 136 500 160
436 141 492 157
7 9V Line
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
823 115 910 139
830 120 902 136
9 3.3V Line
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
